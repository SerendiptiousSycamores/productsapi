CREATE KEYSPACE products WITH replication =
  {‘class’: ‘SimpleStrategy’, ‘replication_factor’ : 1};

/* partition index tells you which node
/* cluster key for sorting
/* can also do a join for related_product

/* query: product info by product id */
CREATE TYPE feature (
  feature text NOT NULL,
  value text NOT NULL
)

CREATE TABLE product (
  productid uuid NOT NULL,
  name text NOT NULL,
  slogan text NOT NULL,
  description text NOT NULL,
  category text NOT NULL,
  default_price int NOT NULL,
  features map<feature> NOT NULL,
  PRIMARY KEY (productid)
);

/* query: find styles by product id */
CREATE TYPE photos (
  url text NOT NULL,
  thumbnail text NOT NULL
)

CREATE TYPE sku (
  size text NOT NULL,
  quantity int NOT NULL
)

CREATE TYPE style (
  name text NOT NULL,
  price int NOT NULL,
  salePrice int NOT NULL,
  default boolean NOT NULL,
  photos map<photos> NOT NULL,
  skus map<text, sku> NOT NULL
)

CREATE TABLE style_by_productid (
  productid int NOT NULL,
  styleid int NOT NULL,
  results map<style> NOT NULL,
  PRIMARY KEY (productid)
);

/* query: find related by product id */
CREATE TABLE related_by_productid (
  productid int NOT NULL,
  relatedid uuid NOT NULL,
  related set<int> NOT NULL,
  PRIMARY KEY (productid)
)

/* query: find skus by style id */
-- CREATE TABLE skus_by_style (
--   styleid int,
--   skuid uuid,
--   sku text,
--   sku map<text, frozen<sku>>,
--   PRIMARY KEY (styleid, skuid),
-- );

-- /* query: find photos by style id */
-- CREATE TYPE photos (
--   url text,
--   thumbnail text
-- )

-- CREATE TABLE photos_by_style (
--   styleid int,
--   photosid uuid,
--   photos map<frozen<photos>>,
--   PRIMARY KEY (styleid, photosid)
-- )

-- psql postgres
-- \CREATE USER <user> WITH PASSWORD <password>;
-- \CREATE ROLE <user> WITH PASSWORD <password>;
-- \ALTER ROLE <user> CREATEDB;
-- psql postgres -U <user>

-- CREATE TABLE skus (
--   id serial,
--   style_id INT,
--   size varchar(5) NOT NULL,
--   quantity INT NOT NULL,
--   PRIMARY KEY (id),
--   FOREIGN KEY (style_id) REFERENCES style (id)
-- );

-- CREATE TABLE photos (
--   id INT AUTO_INCREMENT,
--   style_id INT,
--   url varchar(250) NOT NULL,
--   thumbnail varchar(250) NOT NULL,
--   PRIMARY KEY (id),
--   FOREIGN KEY (style_id) REFERENCES style (id)
-- );


-- /* add features as an array to product */
-- CREATE TABLE features (
--   id serial,
--   product_id INT NOT NUL,
--   feature varchar(50) NOT NULL,
--   value varchar(50) NOT NULL,
--   PRIMARY KEY (id),
--   FOREIGN KEY (product_id) REFERENCES product (id)
-- );

/* psql -U Ika -d products -f schema.sql */

--  default? boolean NOT NULL,